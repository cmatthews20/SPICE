** Profile: "SCHEMATIC1-firstsim"  [ C:\Users\keepi\Downloads\cole4400lab5-PSpiceFiles\SCHEMATIC1\firstsim.sim ] 

** Creating circuit file "firstsim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../cole4400lab5-pspicefiles/cole4400lab5.lib" 
* From [PSPICE NETLIST] section of C:\Users\keepi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 0 15 1 
+ LIN V_V2 0 15 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
